module ex5(x1,x2,x3,x4,f);
input x1, x2, x3, x4;
output f;
//continuous assignment
  assign f=(x1&x2&x4)|(x1&x2&x3)|(x2&x3&x4)|(x1&x3&x4);
endmodule
