module ex1(a,b,c,d,f);
input a, b, c, d;
output f;
//continuous assignment
assign f=((~a)&b)|(c&d)|((~b)&c)|(b&(~c)&(~d));
endmodule
